LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_SIGNED.all;


ENTITY text IS
	PORT
		( clk								: IN std_logic;
        pixel_row, pixel_column	: IN std_logic_vector(9 DOWNTO 0);
		  char_on						: out std_logic);		
END text;

architecture behavior of text is

--Signals for character 1
SIGNAL size 					: std_logic_vector(9 DOWNTO 0) := "0000001111";  
SIGNAL y_pos					: std_logic_vector(9 DOWNTO 0) := "0100110000";
SiGNAL x_pos					: std_logic_vector(9 DOWNTO 0) := "0100110000";
SIGNAL char_A					: std_logic_vector(5 downto 0) := "000001";
SIGNAL char_A_on				: std_logic;         

component char_rom IS
	PORT
	(
		character_address		:	IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		font_row, font_col	:	IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		clock						: 	IN STD_LOGIC ;
		rom_mux_output			:	OUT STD_LOGIC
	);
END component;

BEGIN

--Component for character 1
char_display: char_rom port map(
		character_address => char_A,
		font_row => pixel_row(3 downto 1),
		font_col => pixel_column(3 downto 1),
		clock => clk,
		rom_mux_output => char_A_on);
		

char_on <= 	'1'	when ( ('0' & x_pos <= '0' & pixel_column) and ('0' & pixel_column <= '0' & x_pos + size) 	-- x_pos - size <= pixel_column <= x_pos + size
						and ('0' & y_pos <= pixel_row ) and ('0' & pixel_row <= y_pos + size)	-- y_pos - size <= pixel_row <= y_pos + size
						and (char_A_on = '1')) else
				'0';


END behavior;

